module INSTR_MEM(
    input [4:0] PC,
    output reg [31:0] IR
);

    reg [31:0] INSTR_MEM[0:31]; 

    initial begin
        INSTR_MEM[0]  = 32'b00110100000001000000000000001010; // ori $a0, $0, 10
        INSTR_MEM[1]  = 32'b00110100000001010000000000000001; // ori $a1, $0, 1
        INSTR_MEM[2]  = 32'b00110100000001100000000000000010; // ori $a2, $0, 2
        INSTR_MEM[3]  = 32'b00000000101001100001000000100000; // add $v0, $a1, $a2
        INSTR_MEM[4]  = 32'b00000001100000000010100000100000; // move $a1, $a2
        INSTR_MEM[5]  = 32'b00000000010000000011000000100000; // move $a2, $v0
        INSTR_MEM[6]  = 32'b00100000100001001111111111111111; // addi $a0, $a0, -1
        INSTR_MEM[7]  = 32'b00011100100000001111111111111011; // bgtz $a0, loop
        INSTR_MEM[8]  = 32'b00000000000000000000000000000000; // nop (exit)
        INSTR_MEM[9]  = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[10] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[11] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[12] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[13] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[14] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[15] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[16] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[17] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[18] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[19] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[20] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[21] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[22] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[23] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[24] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[25] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[26] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[27] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[28] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[29] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[30] = 32'b00000000000000000000000000000000; // nop
        INSTR_MEM[31] = 32'b00000000000000000000000000000000; // nop
    end

    always @(PC) begin
        IR = INSTR_MEM[PC];
    end

endmodule
